`timescale 1ns/1ps

module AXITracer #(
    TargetAddrWidth = 64, // max 64
    TargetIDWdith = 4,    // max 128
    TraceAR = 1,
    TraceAW = 1,
    TraceRLast = 1,
    TraceWLast = 1,
    TraceB = 1
) (
    ports
);

endmodule